//! ALU that can perform add, sub, and, or.
//! Additionally output the *ALUOutput is zero* signal to execute branching control.
module ALU(
    input [31:0]    a,  //! rs1
    input [31:0]    b,  //! rs2 / imm
    input [4:0]     ALUCtrl,    //! ALU operation selected from ALU control
    output reg [31:0]   ALUOutput
    //output          ALUBranch
);

//! Select the operation needed based on ALUCtrl, signal generated by ALUControl by decoding instruction.
always@(*) begin : AluOperation
    case(ALUCtrl)
        0: ALUOutput = a + b;                                      //ADD
        1: ALUOutput = a - b;                                      //SUB
        2: ALUOutput = a << b[4:0];                                //SLL
        3: ALUOutput = ($signed(a) < $signed(b)) ? 32'b1 : 32'b0 ; //SLT
        4: ALUOutput = (a < b) ? 32'b1 : 32'b0;                    //SLTU
        5: ALUOutput = a ^ b;                                      //XOR
        6: ALUOutput = a >> b[4:0];                                //SRL  REVISAR QUE FUNCIONEN BIEN
        7: ALUOutput = a >>> b[4:0];                               //SRA  REVISAR QUE FUNCIONEN BIEN
        8: ALUOutput = a | b;                                      //OR
        9: ALUOutput = a & b;                                      //AND
        default: ALUOutput = 0;
    endcase
end

//assign ALUBranch = (ALUOutput==0);

endmodule
